// Deprecated: clock_divider has been renamed to sevenseg_clock_divider.
// This file is intentionally left without a module to prevent duplicate definitions.