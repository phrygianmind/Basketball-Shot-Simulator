`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/26/2025 05:57:56 PM
// Design Name: 
// Module Name: Basketball_Shot
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Basketball_Shot(
    //VGA
    input CLK100MHZ, 
    //input wire reset,             // optional can connect to a button
    output wire [11:0] rgb,
    output wire VGA_HS,
    output wire VGA_VS
    
    //Accelerometer
    
    
    //Seven Seg LED

    );
    
    
    
    
    
    
    
    
    
    
endmodule
